module decay(
    input   wire [0:7]  in,
    output  wire [0:7]  out
);

assign wire 

endmodule