module neuron(
    input   wire [0:8]  inputs,
    input   wire        learn,
    input   wire        clk,
    output  wire        spike_out
);

synapse s0

endmodule